// ============================================================================
// Copyright (c) 2016 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altera Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL/Verilog or C/C++ source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// ============================================================================
//           
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//  
//  
//                     web: http://www.terasic.com/  
//                     email: support@terasic.com
//
// ============================================================================
//Date:  Tue Sep 27 10:46:00 2016
// ============================================================================

`define ENABLE_HPS
`define ENABLE_HSMC

module DE10_Standard_GHRD(


      ///////// CLOCK /////////
      input              CLOCK2_50,
      input              CLOCK3_50,
      input              CLOCK4_50,
      input              CLOCK_50,

      ///////// KEY /////////
      input    [ 3: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LED /////////
      output   [ 9: 0]   LEDR,

      ///////// Seg7 /////////
      output   [ 6: 0]   HEX0,
      output   [ 6: 0]   HEX1,
      output   [ 6: 0]   HEX2,
      output   [ 6: 0]   HEX3,
      output   [ 6: 0]   HEX4,
      output   [ 6: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// Video-In /////////
      input              TD_CLK27,
      input              TD_HS,
      input              TD_VS,
      input    [ 7: 0]   TD_DATA,
      output             TD_RESET_N,

      ///////// VGA /////////
      output             VGA_CLK,
      output             VGA_HS,
      output             VGA_VS,
      output   [ 7: 0]   VGA_R,
      output   [ 7: 0]   VGA_G,
      output   [ 7: 0]   VGA_B,
      output             VGA_BLANK_N,
      output             VGA_SYNC_N,

      ///////// Audio /////////
      inout              AUD_BCLK,
      output             AUD_XCK,
      inout              AUD_ADCLRCK,
      input              AUD_ADCDAT,
      inout              AUD_DACLRCK,
      output             AUD_DACDAT,

      ///////// PS2 /////////
      inout              PS2_CLK,
      inout              PS2_CLK2,
      inout              PS2_DAT,
      inout              PS2_DAT2,

      ///////// ADC /////////
      output             ADC_SCLK,
      input              ADC_DOUT,
      output             ADC_DIN,
      output             ADC_CONVST,

      ///////// I2C for Audio and Video-In /////////
      output             FPGA_I2C_SCLK,
      inout              FPGA_I2C_SDAT,

      ///////// GPIO /////////
      inout    [35: 0]   GPIO,

`ifdef ENABLE_HSMC
      ///////// HSMC /////////
      input              HSMC_CLKIN_P1,
      input              HSMC_CLKIN_N1,
      output             HSMC_CLKIN_P2,
      output             HSMC_CLKIN_N2,
      output             HSMC_CLKOUT_P1,
      output             HSMC_CLKOUT_N1,
      output             HSMC_CLKOUT_P2,
      output             HSMC_CLKOUT_N2,
      inout    [16: 0]   HSMC_TX_D_P,
      inout    [16: 0]   HSMC_TX_D_N,
      inout    [16: 0]   HSMC_RX_D_P,
      inout    [16: 0]   HSMC_RX_D_N,
      input              HSMC_CLKIN0,
      output             HSMC_CLKOUT0,
      inout    [ 3: 0]   HSMC_D,
      output             HSMC_SCL,
      inout              HSMC_SDA,
`endif /*ENABLE_HSMC*/

`ifdef ENABLE_HPS
      ///////// HPS /////////
      inout              HPS_CONV_USB_N,
      output      [14:0] HPS_DDR3_ADDR,
      output      [2:0]  HPS_DDR3_BA,
      output             HPS_DDR3_CAS_N,
      output             HPS_DDR3_CKE,
      output             HPS_DDR3_CK_N,
      output             HPS_DDR3_CK_P,
      output             HPS_DDR3_CS_N,
      output      [3:0]  HPS_DDR3_DM,
      inout       [31:0] HPS_DDR3_DQ,
      inout       [3:0]  HPS_DDR3_DQS_N,
      inout       [3:0]  HPS_DDR3_DQS_P,
      output             HPS_DDR3_ODT,
      output             HPS_DDR3_RAS_N,
      output             HPS_DDR3_RESET_N,
      input              HPS_DDR3_RZQ,
      output             HPS_DDR3_WE_N,
      output             HPS_ENET_GTX_CLK,
      inout              HPS_ENET_INT_N,
      output             HPS_ENET_MDC,
      inout              HPS_ENET_MDIO,
      input              HPS_ENET_RX_CLK,
      input       [3:0]  HPS_ENET_RX_DATA,
      input              HPS_ENET_RX_DV,
      output      [3:0]  HPS_ENET_TX_DATA,
      output             HPS_ENET_TX_EN,
      inout       [3:0]  HPS_FLASH_DATA,
      output             HPS_FLASH_DCLK,
      output             HPS_FLASH_NCSO,
      inout              HPS_GSENSOR_INT,
      inout              HPS_I2C1_SCLK,
      inout              HPS_I2C1_SDAT,
      inout              HPS_I2C2_SCLK,
      inout              HPS_I2C2_SDAT,
      inout              HPS_I2C_CONTROL,
      inout              HPS_KEY,
      inout              HPS_LCM_BK,
      inout              HPS_LCM_D_C,
      inout              HPS_LCM_RST_N,
      output             HPS_LCM_SPIM_CLK,
      output             HPS_LCM_SPIM_MOSI,
      output             HPS_LCM_SPIM_SS,
		input 				 HPS_LCM_SPIM_MISO,
      inout              HPS_LED,
      inout              HPS_LTC_GPIO,
      output             HPS_SD_CLK,
      inout              HPS_SD_CMD,
      inout       [3:0]  HPS_SD_DATA,
      output             HPS_SPIM_CLK,
      input              HPS_SPIM_MISO,
      output             HPS_SPIM_MOSI,
      inout              HPS_SPIM_SS,
      input              HPS_UART_RX,
      output             HPS_UART_TX,
      input              HPS_USB_CLKOUT,
      inout       [7:0]  HPS_USB_DATA,
      input              HPS_USB_DIR,
      input              HPS_USB_NXT,
      output             HPS_USB_STP,
`endif /*ENABLE_HPS*/
      ///////// IR /////////
      output             IRDA_TXD,
      input              IRDA_RXD
);

//=======================================================
//  Fractional PLL START
//=======================================================
	reg fPLL_clock;

	reg [63:0] reconfig_to_pll;
	reg [63:0] reconfig_from_pll;
	reg mgmt_waitrequest;
	reg mgmt_write;
	reg [5:0] mgmt_address;
	reg [31:0] mgmt_writedata;
	
	
	assign LEDR[0] = GPS_signal;

	
	assign HSMC_CLKIN_N2 = fPLL_clock;
	assign HSMC_CLKIN_P2 = GPS_signal;
	
//	assign GPIO[25] = GPS_signal;
//	assign GPIO[21] = fPLL_clock;
//=======================================================
//  Structural coding
//=======================================================
	
	fractional_PLL_1(
		.refclk            (CLOCK_50),            //            refclk.clk
		.rst               (rst),               //             reset.reset
		.outclk_0          (fPLL_clock),          //           outclk0.clk
		.locked            (locked),            //            locked.export
		.reconfig_to_pll   (reconfig_to_pll),   //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (reconfig_from_pll)  // reconfig_from_pll.reconfig_from_pll

	);
	
	
	pll_reconfiguration_1 (
		.mgmt_clk          (CLOCK_50),          //          mgmt_clk.clk
		.mgmt_reset        (mgmt_reset),        //        mgmt_reset.reset
		.mgmt_waitrequest  (mgmt_waitrequest),  // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mgmt_read),         //                  .read
		.mgmt_write        (mgmt_write),        //                  .write
		.mgmt_readdata     (mgmt_readdata),     //                  .readdata
		.mgmt_address      (mgmt_address),      //                  .address
		.mgmt_writedata    (mgmt_writedata),    //                  .writedata
		.reconfig_to_pll   (reconfig_to_pll),   //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (reconfig_from_pll) // reconfig_from_pll.reconfig_from_pll
	);



//=======================================================
//  Structural coding
//=======================================================
	reg [31:0] fPLL_counter = 0;
	reg [31:0] c_out = 0;
	reg [31:0] K_counter = 2147483606 /* synthesis keep */;

	reg [31:0] target = 25000000;
//	wire [31:0] target;
	reg [31:0] error = 0;
	
	reg SM_trig = 0;

	
	
	reg [3:0] fPLL_SM;
	
	wire GPS_signal;
	assign GPS_signal = GPIO[0];
	
	
	always @(posedge fPLL_clock & SW[9])
	begin
		fPLL_counter =  fPLL_counter + 1;
		
		case(SM_trig)
	
			1'b0:
				begin
					if (GPS_signal == 1)
						begin
							if (fPLL_counter < target)
								begin
									c_out = fPLL_counter;
									error = target - fPLL_counter;
									
									if (error > 1000)
										K_counter = K_counter;
									else
										K_counter = K_counter + 5435*error;
										
									fPLL_counter = 0;
									SM_trig = 1'b1;
								end
								
							else if (fPLL_counter > target)
								begin
									c_out = fPLL_counter;
									error = fPLL_counter - target;
									
									if (error > 1000)
										K_counter = K_counter;
									else
										K_counter = K_counter - 5435*error;
	
									fPLL_counter = 0;
									SM_trig = 1'b1;
								end
							else
								begin
									c_out = fPLL_counter;
									error = 0;
									K_counter = K_counter;
									fPLL_counter = 0;
									SM_trig = 1'b1;
								end
						end
				end
				
			1'b1:
				begin
					if (GPS_signal == 0)
						begin
							SM_trig <= 1'b0;
						end
				end
				
		endcase
	
			
		case(fPLL_SM)
		
			4'b0000:
				begin
					if (mgmt_waitrequest == 0 & GPS_signal == 1)
						begin
							mgmt_writedata = 32'd0;
							mgmt_address = 6'b000000;
							fPLL_SM <= 4'b0001;
						end
				end
				
			4'b0001:
				begin
					mgmt_write = 1;
					fPLL_SM <= 4'b0010;
				end
			
			4'b0010:
				begin
					mgmt_write = 0;
					fPLL_SM <= 4'b0011;
				end
				
			4'b0011:
				begin
					mgmt_writedata = K_counter;
					mgmt_address = 6'b000111;
					fPLL_SM <= 4'b0100;
				end
			
			4'b0100:
				begin
					mgmt_write = 1;
					fPLL_SM <= 4'b0101;
				end
				
			4'b0101:
				begin
					mgmt_write = 0;
					fPLL_SM <= 4'b0111;
				end

			4'b0111:
				begin
					mgmt_writedata = 32'd0;
					mgmt_address = 6'b000010;
					fPLL_SM <= 4'b1000;
				end
				
			4'b1000:
				begin
					mgmt_write = 1;
					fPLL_SM <= 4'b1001;
				end
				
			4'b1001:
				begin
					mgmt_write = 0;
					fPLL_SM <= 4'b1011;
				end
				
			4'b1011:
				begin
					if (GPS_signal == 0)
						begin
							fPLL_SM <= 4'b0000;
						end
				end
			
		endcase
	end

//=======================================================
//  Fractional PLL END
//=======================================================




//=======================================================
//  REG/WIRE declarations
//=======================================================

  reg clock_100;
  reg clock_12;
  
  my_pll (
		.refclk   (fPLL_clock),   //  refclk.clk
		.rst      (rst),      //   reset.reset
		.outclk_0 (clock_100), // outclk0.clk
		.outclk_1 (clock_12), // outclk1.clk
		.locked   (locked)    //  locked.export
	);
	
//busybox devmem 0xc5000020 w 0x00000001
//busybox devmem 0xc5000010 w 0x00000001
	
	reg hps_continue = 0;
	reg hps_start = 0;

	assign LEDR[9] = hps_start;

	assign LEDR[1] = GPIO[17];
	assign LEDR[2] = GPIO[5];
	assign LEDR[3] = GPIO[9];
	assign LEDR[4] = GPIO[13];
	
	
//=======================================================
//  Structural coding
//=======================================================
	reg cpy_en_0 = 0;
	reg cpy_en_1 = 0;
	reg cpy_en_2 = 0;
	reg cpy_en_3 = 0;
	
	reg [14:0] addr_0;
	reg [14:0] addr_1;
	reg [14:0] addr_2;
	reg [14:0] addr_3;
	
	reg [31:0] bank_0;
	reg [31:0] bank_1;
	reg [31:0] bank_2;
	reg [31:0] bank_3;
	
	reg [29:0] timetagger;
	
	always @(posedge clock_100 & hps_start)
	begin
		timetagger <= timetagger + 1;
	end
	
////////////////////////////////////////////////////////////	
	always @(posedge r3_Data & hps_start)
	begin
		addr_0 = addr_0 + 1;
		
		if(addr_0 == 16383 | addr_0 == 32767)
			begin
				bank_0 = bank_0 + 1;
				cpy_en_0 = ~cpy_en_0;
			end
	end
	
//////////////////////////////////////////////////////////////	
	
	always @(posedge r6_Data & hps_start)
	begin
		addr_1 = addr_1 + 1;
		
		if(addr_1 == 16383 | addr_1 == 32767)
			begin
				bank_1 = bank_1 + 1;
				cpy_en_1 = ~cpy_en_1;
			end
	end
	
//////////////////////////////////////////////////////////////
	
	always @(posedge r9_Data & hps_start)
	begin
		addr_2 = addr_2 + 1;
		
		if(addr_2 == 16383 | addr_2 == 32767)
			begin
				bank_2 = bank_2 + 1;
				cpy_en_2 = ~cpy_en_2;
			end
	end
	
//////////////////////////////////////////////////////////////
	
	always @(posedge r12_Data & hps_start)
	begin
		addr_3 = addr_3 + 1;
		
		if(addr_3 == 16383 | addr_3 == 32767)
			begin
				bank_3 = bank_3 + 1;
				cpy_en_3 = ~cpy_en_3;
			end
	end
///////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////
	reg r1_Data;
	reg r2_Data;
	reg r3_Data;
	
	reg r4_Data;
	reg r5_Data;
	reg r6_Data;
	
	reg r7_Data;
	reg r8_Data;
	reg r9_Data;
	
	reg r10_Data;
	reg r11_Data;
	reg r12_Data;
	
	
	always @(posedge clock_100)
	begin
	 r1_Data <= GPIO[17];
	 r2_Data <= r1_Data;
	 r3_Data <= r2_Data;
	end
	
	always @(posedge clock_100)
	begin
	 r4_Data <= GPIO[5];
	 r5_Data <= r4_Data;
	 r6_Data <= r5_Data;
	end
	
	always @(posedge clock_100)
	begin
	 r7_Data <= GPIO[9];
	 r8_Data <= r7_Data;
	 r9_Data <= r8_Data;
	end
	
	always @(posedge clock_100)
	begin
	 r10_Data <= GPIO[13];
	 r11_Data <= r10_Data;
	 r12_Data <= r11_Data;
	end
	

//=======================================================
//  REG/WIRE declarations
//=======================================================
  wire  hps_fpga_reset_n;
  wire [3:0] fpga_debounced_buttons;
  wire [8:0]  fpga_led_internal;
  wire [2:0]  hps_reset_req;
  wire        hps_cold_reset;
  wire        hps_warm_reset;
  wire        hps_debug_reset;
  wire [27:0] stm_hw_events;
  wire        fpga_clk_50;
// connection of internal logics
//  assign LEDR[9:1] = fpga_led_internal;
  assign stm_hw_events    = {{4{1'b0}}, SW, fpga_led_internal, fpga_debounced_buttons};
  assign fpga_clk_50=CLOCK_50;
//=======================================================
//  Structural coding
//=======================================================
soc_system u0 (      
		  .clk_clk                               (clock_100),                             //                clk.clk
		  .reset_reset_n                         (1'b1),                                 //                reset.reset_n
		  /////////////////////////////////////////////////////////////////////////////////
		  .mem_0_address                         (addr_0),                              //                     mem_0.address
        .mem_0_chipselect                      (1'b1),                                //                          .chipselect
        .mem_0_clken                           (1'b1),                                 //                          .clken
        .mem_0_write                           (r3_Data & hps_start),                                //                          .write
        .mem_0_readdata                        (),                                     //                          .readdata
        .mem_0_writedata                       (timetagger),                              //                          .writedata
        .mem_0_byteenable                      (4'b1111),                                 //                          .byteenable
		  
		  .mem_1_address                         (addr_1),                              //                     mem_0.address
        .mem_1_chipselect                      (1'b1),                                //                          .chipselect
        .mem_1_clken                           (1'b1),                                 //                          .clken
        .mem_1_write                           (r6_Data & hps_start),                                //                          .write
        .mem_1_readdata                        (),                                     //                          .readdata
        .mem_1_writedata                       (timetagger),                              //                          .writedata
        .mem_1_byteenable                      (4'b1111),                                 //                          .byteenable

		  .mem_2_address                         (addr_2),                              //                     mem_0.address
        .mem_2_chipselect                      (1'b1),                                //                          .chipselect
        .mem_2_clken                           (1'b1),                                 //                          .clken
        .mem_2_write                           (r9_Data & hps_start),                                //                          .write
        .mem_2_readdata                        (),                                     //                          .readdata
        .mem_2_writedata                       (timetagger),                              //                          .writedata
        .mem_2_byteenable                      (4'b1111),                                 //                          .byteenable

		  .mem_3_address                         (addr_3),                              //                     mem_0.address
        .mem_3_chipselect                      (1'b1),                                //                          .chipselect
        .mem_3_clken                           (1'b1),                                 //                          .clken
        .mem_3_write                           (r12_Data & hps_start),                                //                          .write
        .mem_3_readdata                        (),                                     //                          .readdata
        .mem_3_writedata                       (timetagger),                              //                          .writedata
        .mem_3_byteenable                      (4'b1111),                                 //                          .byteenable

		  
		  .adr_count_0_export                    (cpy_en_0),                               //                 adr_count.export
		  .adr_count_1_export                    (cpy_en_1),                               //                 adr_count.export
		  .adr_count_2_export                    (cpy_en_2),                    //               adr_count_2.export
        .adr_count_3_export                    (cpy_en_3),                     //               adr_count_3.export

		  .hps_continue_export                   (hps_continue),                    //              hps_continue.export
		  .hps_start_export                      (hps_start),                       //                 hps_start.export
		  /////////////////////////////////////////////////////////////////////////////////
		  
		  //HPS ddr3
		  .memory_mem_a                          ( HPS_DDR3_ADDR),                       //                memory.mem_a
        .memory_mem_ba                         ( HPS_DDR3_BA),                         //                .mem_ba
        .memory_mem_ck                         ( HPS_DDR3_CK_P),                       //                .mem_ck
        .memory_mem_ck_n                       ( HPS_DDR3_CK_N),                       //                .mem_ck_n
        .memory_mem_cke                        ( HPS_DDR3_CKE),                        //                .mem_cke
        .memory_mem_cs_n                       ( HPS_DDR3_CS_N),                       //                .mem_cs_n
        .memory_mem_ras_n                      ( HPS_DDR3_RAS_N),                      //                .mem_ras_n
        .memory_mem_cas_n                      ( HPS_DDR3_CAS_N),                      //                .mem_cas_n
        .memory_mem_we_n                       ( HPS_DDR3_WE_N),                       //                .mem_we_n
        .memory_mem_reset_n                    ( HPS_DDR3_RESET_N),                    //                .mem_reset_n
        .memory_mem_dq                         ( HPS_DDR3_DQ),                         //                .mem_dq
        .memory_mem_dqs                        ( HPS_DDR3_DQS_P),                      //                .mem_dqs
        .memory_mem_dqs_n                      ( HPS_DDR3_DQS_N),                      //                .mem_dqs_n
        .memory_mem_odt                        ( HPS_DDR3_ODT),                        //                .mem_odt
        .memory_mem_dm                         ( HPS_DDR3_DM),                         //                .mem_dm
        .memory_oct_rzqin                      ( HPS_DDR3_RZQ),                        //                .oct_rzqin
       //HPS ethernet		
	     .hps_0_hps_io_hps_io_emac1_inst_TX_CLK ( HPS_ENET_GTX_CLK),       //                             hps_0_hps_io.hps_io_emac1_inst_TX_CLK
        .hps_0_hps_io_hps_io_emac1_inst_TXD0   ( HPS_ENET_TX_DATA[0] ),   //                             .hps_io_emac1_inst_TXD0
        .hps_0_hps_io_hps_io_emac1_inst_TXD1   ( HPS_ENET_TX_DATA[1] ),   //                             .hps_io_emac1_inst_TXD1
        .hps_0_hps_io_hps_io_emac1_inst_TXD2   ( HPS_ENET_TX_DATA[2] ),   //                             .hps_io_emac1_inst_TXD2
        .hps_0_hps_io_hps_io_emac1_inst_TXD3   ( HPS_ENET_TX_DATA[3] ),   //                             .hps_io_emac1_inst_TXD3
        .hps_0_hps_io_hps_io_emac1_inst_RXD0   ( HPS_ENET_RX_DATA[0] ),   //                             .hps_io_emac1_inst_RXD0
        .hps_0_hps_io_hps_io_emac1_inst_MDIO   ( HPS_ENET_MDIO ),         //                             .hps_io_emac1_inst_MDIO
        .hps_0_hps_io_hps_io_emac1_inst_MDC    ( HPS_ENET_MDC  ),         //                             .hps_io_emac1_inst_MDC
        .hps_0_hps_io_hps_io_emac1_inst_RX_CTL ( HPS_ENET_RX_DV),         //                             .hps_io_emac1_inst_RX_CTL
        .hps_0_hps_io_hps_io_emac1_inst_TX_CTL ( HPS_ENET_TX_EN),         //                             .hps_io_emac1_inst_TX_CTL
        .hps_0_hps_io_hps_io_emac1_inst_RX_CLK ( HPS_ENET_RX_CLK),        //                             .hps_io_emac1_inst_RX_CLK
        .hps_0_hps_io_hps_io_emac1_inst_RXD1   ( HPS_ENET_RX_DATA[1] ),   //                             .hps_io_emac1_inst_RXD1
        .hps_0_hps_io_hps_io_emac1_inst_RXD2   ( HPS_ENET_RX_DATA[2] ),   //                             .hps_io_emac1_inst_RXD2
        .hps_0_hps_io_hps_io_emac1_inst_RXD3   ( HPS_ENET_RX_DATA[3] ),   //                             .hps_io_emac1_inst_RXD3
       //HPS QSPI  
		  .hps_0_hps_io_hps_io_qspi_inst_IO0     ( HPS_FLASH_DATA[0]    ),     //                               .hps_io_qspi_inst_IO0
        .hps_0_hps_io_hps_io_qspi_inst_IO1     ( HPS_FLASH_DATA[1]    ),     //                               .hps_io_qspi_inst_IO1
        .hps_0_hps_io_hps_io_qspi_inst_IO2     ( HPS_FLASH_DATA[2]    ),     //                               .hps_io_qspi_inst_IO2
        .hps_0_hps_io_hps_io_qspi_inst_IO3     ( HPS_FLASH_DATA[3]    ),     //                               .hps_io_qspi_inst_IO3
        .hps_0_hps_io_hps_io_qspi_inst_SS0     ( HPS_FLASH_NCSO    ),        //                               .hps_io_qspi_inst_SS0
        .hps_0_hps_io_hps_io_qspi_inst_CLK     ( HPS_FLASH_DCLK    ),        //                               .hps_io_qspi_inst_CLK
       //HPS SD card 
		  .hps_0_hps_io_hps_io_sdio_inst_CMD     ( HPS_SD_CMD    ),           //                               .hps_io_sdio_inst_CMD
        .hps_0_hps_io_hps_io_sdio_inst_D0      ( HPS_SD_DATA[0]     ),      //                               .hps_io_sdio_inst_D0
        .hps_0_hps_io_hps_io_sdio_inst_D1      ( HPS_SD_DATA[1]     ),      //                               .hps_io_sdio_inst_D1
        .hps_0_hps_io_hps_io_sdio_inst_CLK     ( HPS_SD_CLK   ),            //                               .hps_io_sdio_inst_CLK
        .hps_0_hps_io_hps_io_sdio_inst_D2      ( HPS_SD_DATA[2]     ),      //                               .hps_io_sdio_inst_D2
        .hps_0_hps_io_hps_io_sdio_inst_D3      ( HPS_SD_DATA[3]     ),      //                               .hps_io_sdio_inst_D3
       //HPS USB 		  
		  .hps_0_hps_io_hps_io_usb1_inst_D0      ( HPS_USB_DATA[0]    ),      //                               .hps_io_usb1_inst_D0
        .hps_0_hps_io_hps_io_usb1_inst_D1      ( HPS_USB_DATA[1]    ),      //                               .hps_io_usb1_inst_D1
        .hps_0_hps_io_hps_io_usb1_inst_D2      ( HPS_USB_DATA[2]    ),      //                               .hps_io_usb1_inst_D2
        .hps_0_hps_io_hps_io_usb1_inst_D3      ( HPS_USB_DATA[3]    ),      //                               .hps_io_usb1_inst_D3
        .hps_0_hps_io_hps_io_usb1_inst_D4      ( HPS_USB_DATA[4]    ),      //                               .hps_io_usb1_inst_D4
        .hps_0_hps_io_hps_io_usb1_inst_D5      ( HPS_USB_DATA[5]    ),      //                               .hps_io_usb1_inst_D5
        .hps_0_hps_io_hps_io_usb1_inst_D6      ( HPS_USB_DATA[6]    ),      //                               .hps_io_usb1_inst_D6
        .hps_0_hps_io_hps_io_usb1_inst_D7      ( HPS_USB_DATA[7]    ),      //                               .hps_io_usb1_inst_D7
        .hps_0_hps_io_hps_io_usb1_inst_CLK     ( HPS_USB_CLKOUT    ),       //                               .hps_io_usb1_inst_CLK
        .hps_0_hps_io_hps_io_usb1_inst_STP     ( HPS_USB_STP    ),          //                               .hps_io_usb1_inst_STP
        .hps_0_hps_io_hps_io_usb1_inst_DIR     ( HPS_USB_DIR    ),          //                               .hps_io_usb1_inst_DIR
        .hps_0_hps_io_hps_io_usb1_inst_NXT     ( HPS_USB_NXT    ),          //                               .hps_io_usb1_inst_NXT
		  
		  //HPS SPI0->LCDM 	
        .hps_0_hps_io_hps_io_spim0_inst_CLK    ( HPS_LCM_SPIM_CLK),    //                               .hps_io_spim0_inst_CLK
        .hps_0_hps_io_hps_io_spim0_inst_MOSI   ( HPS_LCM_SPIM_MOSI),   //                               .hps_io_spim0_inst_MOSI
        .hps_0_hps_io_hps_io_spim0_inst_MISO   ( HPS_LCM_SPIM_MISO),   //                               .hps_io_spim0_inst_MISO
        .hps_0_hps_io_hps_io_spim0_inst_SS0    ( HPS_LCM_SPIM_SS),    //                               .hps_io_spim0_inst_SS0
       //HPS SPI1 		  
		  .hps_0_hps_io_hps_io_spim1_inst_CLK    ( HPS_SPIM_CLK  ),           //                               .hps_io_spim1_inst_CLK
        .hps_0_hps_io_hps_io_spim1_inst_MOSI   ( HPS_SPIM_MOSI ),           //                               .hps_io_spim1_inst_MOSI
        .hps_0_hps_io_hps_io_spim1_inst_MISO   ( HPS_SPIM_MISO ),           //                               .hps_io_spim1_inst_MISO
        .hps_0_hps_io_hps_io_spim1_inst_SS0    ( HPS_SPIM_SS ),             //                               .hps_io_spim1_inst_SS0
      //HPS UART		
		  .hps_0_hps_io_hps_io_uart0_inst_RX     ( HPS_UART_RX    ),          //                               .hps_io_uart0_inst_RX
        .hps_0_hps_io_hps_io_uart0_inst_TX     ( HPS_UART_TX    ),          //                               .hps_io_uart0_inst_TX
		//HPS I2C1
		  .hps_0_hps_io_hps_io_i2c0_inst_SDA     ( HPS_I2C1_SDAT    ),        //                               .hps_io_i2c0_inst_SDA
        .hps_0_hps_io_hps_io_i2c0_inst_SCL     ( HPS_I2C1_SCLK    ),        //                               .hps_io_i2c0_inst_SCL
		//HPS I2C2
		  .hps_0_hps_io_hps_io_i2c1_inst_SDA     ( HPS_I2C2_SDAT    ),        //                               .hps_io_i2c1_inst_SDA
        .hps_0_hps_io_hps_io_i2c1_inst_SCL     ( HPS_I2C2_SCLK    ),        //                               .hps_io_i2c1_inst_SCL
      //HPS GPIO  
		  .hps_0_hps_io_hps_io_gpio_inst_GPIO09  ( HPS_CONV_USB_N),           //                               .hps_io_gpio_inst_GPIO09
        .hps_0_hps_io_hps_io_gpio_inst_GPIO35  ( HPS_ENET_INT_N),           //                               .hps_io_gpio_inst_GPIO35
        .hps_0_hps_io_hps_io_gpio_inst_GPIO37  ( HPS_LCM_BK ),  //                               .hps_io_gpio_inst_GPIO37
		  .hps_0_hps_io_hps_io_gpio_inst_GPIO40  ( HPS_LTC_GPIO ),              //                               .hps_io_gpio_inst_GPIO40
        .hps_0_hps_io_hps_io_gpio_inst_GPIO41  ( HPS_LCM_D_C ),              //                               .hps_io_gpio_inst_GPIO41
        .hps_0_hps_io_hps_io_gpio_inst_GPIO44  ( HPS_LCM_RST_N  ),  //                               .hps_io_gpio_inst_GPIO44
		  .hps_0_hps_io_hps_io_gpio_inst_GPIO48  ( HPS_I2C_CONTROL),          //                               .hps_io_gpio_inst_GPIO48
        .hps_0_hps_io_hps_io_gpio_inst_GPIO53  ( HPS_LED),                  //                               .hps_io_gpio_inst_GPIO53
        .hps_0_hps_io_hps_io_gpio_inst_GPIO54  ( HPS_KEY),                  //                               .hps_io_gpio_inst_GPIO54
    	  .hps_0_hps_io_hps_io_gpio_inst_GPIO61  ( HPS_GSENSOR_INT),  //                               .hps_io_gpio_inst_GPIO61

			
		  .hps_0_h2f_reset_reset_n               ( hps_fpga_reset_n ),                //                hps_0_h2f_reset.reset_n
		  .hps_0_f2h_cold_reset_req_reset_n      (~hps_cold_reset ),      //       hps_0_f2h_cold_reset_req.reset_n
		  .hps_0_f2h_debug_reset_req_reset_n     (~hps_debug_reset ),     //      hps_0_f2h_debug_reset_req.reset_n
		  .hps_0_f2h_stm_hw_events_stm_hwevents  (stm_hw_events ),  //        hps_0_f2h_stm_hw_events.stm_hwevents
		  .hps_0_f2h_warm_reset_req_reset_n      (~hps_warm_reset ),      //       hps_0_f2h_warm_reset_req.reset_n
  
    );

	 
	 // Debounce logic to clean out glitches within 1ms
debounce debounce_inst (
  .clk                                  (fpga_clk_50),
  .reset_n                              (hps_fpga_reset_n),  
  .data_in                              (KEY),
  .data_out                             (fpga_debounced_buttons)
);
  defparam debounce_inst.WIDTH = 4;
  defparam debounce_inst.POLARITY = "LOW";
  defparam debounce_inst.TIMEOUT = 50000;               // at 50Mhz this is a debounce time of 1ms
  defparam debounce_inst.TIMEOUT_WIDTH = 16;            // ceil(log2(TIMEOUT))
  
// Source/Probe megawizard instance
hps_reset hps_reset_inst (
  .source_clk (fpga_clk_50),
  .source     (hps_reset_req)
);

altera_edge_detector pulse_cold_reset (
  .clk       (fpga_clk_50),
  .rst_n     (hps_fpga_reset_n),
  .signal_in (hps_reset_req[0]),
  .pulse_out (hps_cold_reset)
);
  defparam pulse_cold_reset.PULSE_EXT = 6;
  defparam pulse_cold_reset.EDGE_TYPE = 1;
  defparam pulse_cold_reset.IGNORE_RST_WHILE_BUSY = 1;

altera_edge_detector pulse_warm_reset (
  .clk       (fpga_clk_50),
  .rst_n     (hps_fpga_reset_n),
  .signal_in (hps_reset_req[1]),
  .pulse_out (hps_warm_reset)
);
  defparam pulse_warm_reset.PULSE_EXT = 2;
  defparam pulse_warm_reset.EDGE_TYPE = 1;
  defparam pulse_warm_reset.IGNORE_RST_WHILE_BUSY = 1;
  
altera_edge_detector pulse_debug_reset (
  .clk       (fpga_clk_50),
  .rst_n     (hps_fpga_reset_n),
  .signal_in (hps_reset_req[2]),
  .pulse_out (hps_debug_reset)
);
  defparam pulse_debug_reset.PULSE_EXT = 32;
  defparam pulse_debug_reset.EDGE_TYPE = 1;
  defparam pulse_debug_reset.IGNORE_RST_WHILE_BUSY = 1;
  
reg [25:0] counter; 
reg  led_level;
always @(posedge fpga_clk_50 or negedge hps_fpga_reset_n)
begin
if(~hps_fpga_reset_n)
begin
                counter<=0;
                led_level<=0;
end

else if(counter==24999999)
        begin
                counter<=0;
                led_level<=~led_level;
        end
else
                counter<=counter+1'b1;
end

//assign LEDR[0]=led_level;
endmodule

  